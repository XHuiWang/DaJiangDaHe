`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 

// Author: XHuiWang
//////////////////////////////////////////////////////////////////////////////////


//1024项，存过去两次的跳转情况，初始化为00，表示过去两次均不跳转

// module BHR(
//     //
//     input  clk,
//     input  rstn,
//     //预测端
//     input  [31:0] pc,
//     output logic [1:0]  bhr,
//     //更新端
//     input  update,
//     input  [31:0] update_pc,

//     );
// endmodule
