// -*- Verilog -*-

//`ifdef VERILATOR
`define DIFFTEST_EN
// `define CLAP_CONFIG_BR_PROFILE
// `define CLAP_CONFIG_INST_PROFILE
// `define CLAP_CONFIG_AXI_PROFILE
// `define CLAP_CONFIG_LD_ST_PROFILE
// `define CLAP_CONFIG_CACHE_PROFILE
//`endif
