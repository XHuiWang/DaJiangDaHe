`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/07/21 20:26:04
// Design Name: 
// Module Name: br_pre_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// Author: XHuiWang
//////////////////////////////////////////////////////////////////////////////////


module br_pre_top(

    );
endmodule
